library IEEE;
use IEEE.Std_Logic_1164.all;

entity UART-IP-CORE-VHDL is

end UART-IP-CORE-VHDL;

architecture BEHAV of UART-IP-CORE-VHDL is
--	BEGIN Signals declaration	--


--	END Signals declaration		--
begin 
--Concurrential

end BEHAV;